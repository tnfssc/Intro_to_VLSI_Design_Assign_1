.title Problem 2.1

Vin v1 gnd dc=2.5
R1 v1 v2 2k
VB1 v2 v3 dc=0.7 
R2 v3 v4 2k
VB2 v4 gnd dc=0.7

.control
op
print i(Vin)
.endc
.end
