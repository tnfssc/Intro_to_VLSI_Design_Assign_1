.title Problem 1.1

Vin gnd v1 2.5v
R1 v1 v2 1k
C1 v2 v3 1u
R_s v3 gnd 100
.op

.control
run
print v(v2)
exit
.endc
.end
